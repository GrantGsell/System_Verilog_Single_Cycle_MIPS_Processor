`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Grant Gsell
// 
// Create Date: 11/24/2019 11:24:32 PM
// Module Name: tb_overall_simulation
// Project Name: CPU_Design
//////////////////////////////////////////////////////////////////////////////////
module tb_overall_simulation();
    //Mux Testbecnh
    //tb_mux_2x1 u0();
    //Adder Testbench
    //tb_full_adder_one_bit u1();
    //tb_full_adder_four_bit u2();
    //tb_full_adder_sixteen_bit u3();
    //tb_full_adder_thirtytwo_bit u4();

endmodule
