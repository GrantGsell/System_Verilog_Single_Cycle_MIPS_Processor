`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Grant Gsell 
// 
// Create Date: 11/27/2019 12:50:55 PM
// Module Name: instruction_memory
// Project Name: CPU_Design
//////////////////////////////////////////////////////////////////////////////////
module instruction_memory(
    output [31:0] instruction,
    input [31:0] read_Addr_From_PC,
    input rst
    );
        
    //Internal Signal Instantiations
    logic [31:0] rom [31:0];
    logic [5:0] shifted_Addr;
    
    //Synchronous Block
    always @(posedge rst) begin
        for(integer i=0; i<32; i++) begin
            rom[i] = 32'b0;
        end

        //Test Equation Program
        rom[0] = {6'b001000, 5'b00000, 5'b00001, 16'd1000};                     //addi r1, r0, 1000
        rom[1] = {6'b001000, 5'b00000, 5'b00010, 16'd200};                      //addi r2, r0, 200
        rom[2] = {6'b001000, 5'b00000, 5'b00011, -16'd300};                     //addi r3, r0, -300
        rom[3] = {6'b001000, 5'b00000, 5'b00100, 16'd400};                      //addi r4, r0, 400
        rom[4] = {6'b001000, 5'b00000, 5'b00101, -16'd100};                     //addi r5, r0, -100
        rom[5] = {6'b001000, 5'b00000, 5'b00110, 16'd3};                        //addi r6, r0, 3
        rom[6] = {6'b101011, 5'b00000, 5'b00001, 16'd0};                        //sw r1, 0(0)
        rom[7] = {6'b101011, 5'b00000, 5'b00010, 16'd4};                        //sw r2, 4(0)
        rom[8] = {6'b101011, 5'b00000, 5'b00011, 16'd8};                        //sw r3, 8(0)
        rom[9] = {6'b101011, 5'b00000, 5'b00100, 16'd12};                       //sw r4, 12(0)
        rom[10] = {6'b101011, 5'b00000, 5'b00101, 16'd16};                      //sw r5, 16(0)
        rom[11] = {6'b101011, 5'b00000, 5'b00110, 16'd20};                      //sw r6, 20(0)
        rom[12] = {6'b100011, 5'b00000, 5'b00111, 16'd0};                       //lw r7, 0(0)
        rom[13] = {6'b100011, 5'b00000, 5'b01000, 16'd4};                       //lw r8, 4(0)
        rom[14] = {6'b100011, 5'b00000, 5'b01001, 16'd8};                       //lw r9, 8(0)
        rom[15] = {6'b100011, 5'b00000, 5'b01010, 16'd12};                      //lw r10, 12(0)
        rom[16] = {6'b100011, 5'b00000, 5'b01011, 16'd16};                      //lw r11, 16(0)
        rom[17] = {6'b100011, 5'b00000, 5'b01100, 16'd20};                      //lw r12, 20(0)
        rom[18] = {6'b000000, 5'b00111, 5'b01000, 5'b00111, 11'b00000010010};   //mult r7, r7, r8
        rom[19] = {6'b000000, 5'b01001, 5'b01010, 5'b01001, 11'b00000010010};   //mult r9, r9, r10
        rom[20] = {6'b000000, 5'b00111, 5'b01001, 5'b00111, 11'b00000100000};   //add r7, r7, r9
        rom[21] = {6'b000000, 5'b00111, 5'b01011, 5'b00111, 11'b00000100010};   //sub r7, r7, r11
        rom[22] = {6'b000000, 5'b00111, 5'b01100, 5'b00111, 11'b00000011010};   //div r7, r7, r12
        rom[23] = {6'b101011, 5'b00000, 5'b00111, 16'd28};                      //sw r7, 28(0)
        
        /*
        //Instruction Set Validity Test
        rom[0] = {6'b001000, 5'b00000, 5'b00001, 16'd100};                      //addi r1, r0, 100
        rom[1] = {6'b001000, 5'b00000, 5'b00010, 16'd1};                        //addi r2, r0, 1
        rom[2] = {6'b000000, 5'b00010, 5'b00001, 5'b00011, 11'b00000100000};    //add r3, r2, r1
        rom[3] = {6'b000000, 5'b00011, 5'b00010, 5'b00011, 11'b00000100010};    //sub r3, r3, r2
        rom[4] = {6'b001000, 5'b00000, 5'b00100, 16'd2};                        //addi r4, r0, 2
        rom[5] = {6'b000000, 5'b00011, 5'b00100, 5'b00011, 11'b00000011010};    //div r3, r3, r4
        rom[6] = {6'b000000, 5'b00100, 5'b00010, 5'b00100, 11'b00000100000};    //add r4, r4, r2
        rom[7] = {6'b000000, 5'b00011, 5'b00100, 5'b00011, 11'b00000010010};    //mult r3, r3, r4
        rom[8] = {6'b001000, 5'b00000, 5'b00010, 16'd6};                        //addi r2, r0, 6
        rom[9] = {6'b000000, 5'b00010, 5'b00011, 5'b00011, 11'b00000101000};    //and r3, r3, r2
        rom[10] = {6'b000000, 5'b00001, 5'b00011, 5'b00011, 11'b00000100101};   //or r3, r3, r1
        rom[11] = {6'b001000, 5'b00000, 5'b00010, 16'd9};                       //addi r2, r0, 9
        rom[12] = {6'b000000, 5'b00010, 5'b00011, 5'b00011, 11'b00000100110};   //xor r3, r3, r2
        rom[13] = {6'b101011, 5'b00000, 5'b00011, 16'd0};                       //sw r3, 0(0)
        rom[14] = {6'b101011, 5'b00000, 5'b00010, 16'd4};                       //sw r2, 4(0)
        rom[15] = {6'b100011, 5'b00000, 5'b00110, 16'd0};                       //lw r6, 0(1)
        rom[16] = {6'b100011, 5'b00000, 5'b00101, 16'd4};                       //lw r5, 4(0)
        rom[17] = {6'b001000, 5'b00000, 5'b00111, 16'd115};                     //addi r7, r0, 115
        rom[18] = {6'b001000, 5'b00110, 5'b00110, 16'd4};                       //addi r6, r6, 4
        rom[19] = {6'b000100, 5'b00111, 5'b00110, -16'd2};                      //beq r7, r6, pcAddr-8 (returns to ROM 18)
        rom[20] = {6'b000010, 26'd0};                                           //Jump rom[0]
        */
    end

    assign shifted_Addr = read_Addr_From_PC[6:2];
    assign instruction = rom[shifted_Addr];
endmodule
