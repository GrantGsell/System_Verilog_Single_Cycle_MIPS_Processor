`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Engineer: Grant Gsell
// 
// Create Date: 11/29/2019 09:33:17 PM
// Module Name: tb_instruction_memory
// Project Name: CPU_Design
//////////////////////////////////////////////////////////////////////////////////
module tb_instruction_memory();

endmodule
